//Subject:     CO project 2 - Decoder
//--------------------------------------------------------------------------------
//Version:     1
//--------------------------------------------------------------------------------
//Writer:      Luke
//----------------------------------------------
//Date:        2010/8/16
//----------------------------------------------
//Description: 
//--------------------------------------------------------------------------------

module Decoder(
    instr_op_i,
	RegWrite_o,
	ALU_op_o,
	ALUSrc_o,
	RegDst_o,
	Branch_o,
	//***************************************************
	BranchType_o,
	Jump_o,
	MemRead_o,
	MemWrite_o,
	MemtoReg_o
	);
     
//I/O ports
input  [6-1:0] instr_op_i;

output         RegWrite_o;
output [3-1:0] ALU_op_o;
output [1:0]   ALUSrc_o;
output         RegDst_o;
output         Branch_o;
output	BranchType_o,
output	Jump_o,
output	MemRead_o,
output	MemWrite_o,
output	MemtoReg_o
 
//Internal Signals
reg    [3-1:0] ALU_op_o;
reg    [1:0]   ALUSrc_o;
reg            RegWrite_o;
reg            RegDst_o;
reg            Branch_o;

//Parameter


//Main function
always@(*)begin
	case(instr_op_i)
		6'b000000:begin			//R-type
			ALU_op_o <= 3'b010;
            ALUSrc_o <= 2'b00;
            RegWrite_o <= 1;
            RegDst_o <= 1;
            Branch_o <= 0;
			//FIX ME Here! what is the branchType 
			BranchType_o <=0;     
			Jump_o <= 0;
			MemRead_o <= 0;
			MemWrite_o <= 0;
			MemtoReg_o	<= 0;		
		end
		6'b001000:begin			//ADDI			
			ALU_op_o <= 3'b100;
            ALUSrc_o <= 2'b01;
            RegWrite_o <= 1;
            RegDst_o <= 0;
            Branch_o <= 0;	
			//FIX ME Here! what is the branchType 
			BranchType_o <=0;     
			Jump_o <= 0;
			MemRead_o <= 0;
			MemWrite_o <= 0;
			MemtoReg_o	<= 0;		
		end
		6'b001101:begin			//ORI
		    ALU_op_o <= 3'b101;
            ALUSrc_o <= 2'b10;
            RegWrite_o <= 1;
            RegDst_o <= 0;
            Branch_o <= 0;
			//FIX ME Here! what is the branchType 
			BranchType_o <=0;     
			Jump_o <= 0;
			MemRead_o <= 0;
			MemWrite_o <= 0;
			MemtoReg_o	<= 0;		
		end
		6'b000100:begin			//BEQ
		    ALU_op_o <= 3'b001;
            ALUSrc_o <= 2'b00;
            RegWrite_o <= 0;
            RegDst_o <= 0;		//or X
            Branch_o <= 1;			
			//FIX ME Here! what is the branchType 
			BranchType_o <=0;     
			Jump_o <= 0;
			MemRead_o <= 0;
			MemWrite_o <= 0;
			MemtoReg_o	<= 0;		
		end
		6'b100011:begin			//lw
		    ALU_op_o <= 3'b000;
            ALUSrc_o <= 2'b01;
            RegWrite_o <= 1;
            RegDst_o <= 0;		
            Branch_o <= 0;			
			//FIX ME Here! what is the branchType 
			BranchType_o <=0;     
			Jump_o <= 0;
			MemRead_o <= 1;
			MemWrite_o <= 0;
			MemtoReg_o	<= 1;		
		end		
		6'b101011:begin			//sw
		    ALU_op_o <= 3'b000;
            ALUSrc_o <= 2'b01;
            RegWrite_o <= 0;
            RegDst_o <= 0;		//or X
            Branch_o <= 0;			
			//FIX ME Here! what is the branchType 
			BranchType_o <=0;     
			Jump_o <= 0;
			MemRead_o <= 0;
			MemWrite_o <= 1;
			MemtoReg_o	<= 0;    //or X		
		end
		6'b000010:begin			//jump
		    ALU_op_o <= 3'b000;	//or X
            ALUSrc_o <= 2'b00;	//or X
            RegWrite_o <= 0;	
            RegDst_o <= 0;		//or X
            Branch_o <= 0;			
			//FIX ME Here! what is the branchType 
			BranchType_o <=0;     
			Jump_o <= 1;
			MemRead_o <= 0;
			MemWrite_o <= 0;
			MemtoReg_o	<= 0;    		
		end
	endcase
end

endmodule





                    
                    